LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY decodificador_1a2 IS
	PORT(	w	:IN STD_LOGIC;
			En	:IN STD_LOGIC;
			y	:OUT STD_LOGIC_VECTOR(1 DOWNTO 0));
END decodificador_1a2;

ARCHITECTURE Behavior of decodificador_1a2 IS
	SIGNAL Enw: STD_LOGIC_VECTOR(1 DOWNTO 0);
BEGIN
	Enw <=En&w;
	WITH Enw SELECT
		y<="01" WHEN "10",
			"10" WHEN "11",
			"00" WHEN OTHERS;
END Behavior;