LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY decodificador_columna_verde IS
	PORT(	w	:IN STD_LOGIC_VECTOR(5 DOWNTO 0);
			En	:IN STD_LOGIC;
			y	:OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END decodificador_columna_verde;

ARCHITECTURE Behavior of decodificador_columna_verde IS
	SIGNAL Enw: STD_LOGIC_VECTOR(6 DOWNTO 0);
BEGIN
	Enw <=En&w;
	WITH Enw SELECT
		y<="1111" WHEN "1000000",
			"1110" WHEN "1000001",
			"1110" WHEN "1000010",
			"1110" WHEN "1000011",
			"1110" WHEN "1000100",
			"1110" WHEN "1000101",
			"1110" WHEN "1000110",
			"1110" WHEN "1000111",
			"1110" WHEN "1001000",
			"1100" WHEN "1001001",
			"1100" WHEN "1001010",
			"1100" WHEN "1001011",
			"1100" WHEN "1001100",
			"1100" WHEN "1001101",
			"1100" WHEN "1001110",
			"1100" WHEN "1001111",
			"1100" WHEN "1010000",
			"1000" WHEN "1010001",
			"1000" WHEN "1010010",
			"1000" WHEN "1010011",
			"1000" WHEN "1010100",
			"1000" WHEN "1010101",
			"1000" WHEN "1010110",
			"1000" WHEN "1010111",
			"1000" WHEN "1011000",
			"0000" WHEN "1011001",
			"0000" WHEN "1011010",
			"0000" WHEN "1011011",
			"0000" WHEN "1011100",
			"0000" WHEN "1011101",
			"0000" WHEN "1011110",
			"0000" WHEN "1011111",
			"0000" WHEN "1100000",
			"0000" WHEN "1100001",
			"0000" WHEN "1100010",
			"0000" WHEN "1100011",
			"0000" WHEN "1100100",
			"0000" WHEN "1100101",
			"0000" WHEN "1100110",
			
			"1111" WHEN OTHERS;
END Behavior;