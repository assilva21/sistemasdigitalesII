LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY decodificador_matriz4 IS
	PORT(	w	:IN STD_LOGIC_VECTOR(5 DOWNTO 0);
			En	:IN STD_LOGIC;
			y	:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END decodificador_matriz4;

ARCHITECTURE Behavior of decodificador_matriz4 IS
	SIGNAL Enw: STD_LOGIC_VECTOR(6 DOWNTO 0);
BEGIN
	Enw <=En&w;
	WITH Enw SELECT
		y<="00000000" WHEN "1000000",
			"00000000" WHEN "1000001",
			"00000000" WHEN "1000010",
			"00000000" WHEN "1000011",
			"00000000" WHEN "1000100",
			"00000000" WHEN "1000101",
			"00000000" WHEN "1000110",
			"00000000" WHEN "1000111",
			"00000000" WHEN "1001000",
			"00000000" WHEN "1001001",
			"00000000" WHEN "1001010",
			"00000000" WHEN "1001011",
			"00000000" WHEN "1001100",
			"00000000" WHEN "1001101",
			"00000000" WHEN "1001110",
			"00000000" WHEN "1001111",
			"00000000" WHEN "1010000",
			"00000000" WHEN "1010001",
			"00000000" WHEN "1010010",
			"00000000" WHEN "1010011",
			"00000000" WHEN "1010100",
			"00000000" WHEN "1010101",
			"00000000" WHEN "1010110",
			"00000000" WHEN "1010111",
			"00000000" WHEN "1011000",
			"10000000" WHEN "1011001",
			"11000000" WHEN "1011010",
			"11100000" WHEN "1011011",
			"11110000" WHEN "1011100",
			"11111000" WHEN "1011101",
			"11111100" WHEN "1011110",
			"11111110" WHEN "1011111",
			"11111111" WHEN "1100000",
			"11111111" WHEN "1100001",
			"11111111" WHEN "1100010",
			"11111111" WHEN "1100011",
			"11111111" WHEN "1100100",
			"11111111" WHEN "1100101",
			"11111111" WHEN "1100110",
			"00000000" WHEN OTHERS;
END Behavior;